`ifndef _MY_CONSTANTS_VH_
`define _MY_CONSTANTS_VH_

`timescale 1ns/1ps
`define DUMP_FILE "simulation/waveform.vcd"

`endif // _MY_CONSTANTS_VH_